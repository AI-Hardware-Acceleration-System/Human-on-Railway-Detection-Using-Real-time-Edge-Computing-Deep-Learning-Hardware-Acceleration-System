module FC_tb();
     
parameter datawidth = 16;
parameter input_nodes = 784;
parameter output_nodes = 2;
parameter Mult_Add_Units = 16;

reg clk, reset;
reg [3:0] state;
reg [datawidth*Mult_Add_Units-1:0] input_data;

wire [datawidth*output_nodes-1:0] output_data;
wire done;

Fully_Connect FC(clk,reset,state,input_data,output_data, done);

initial begin
    clk = 0;
    reset = 1;
    state = 1;
    input_data <= 0;
    #15 reset = 0;
    #10 reset = 1;
    state = 11;
    #10 input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10 input_data = 256'h4200_4200_4200_4200_4200_4200_4200_42004200_4200_4200_42004200_4200_4200_4200;
    #10 input_data = 256'h4400_4400_4400_44004400_4400_4400_44004400_4400_4400_44004400_4400_4400_4400;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h0;
    #30input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 256'h4000_4000_4000_4000_4000_4000_4000_40004000_4000_4000_40004000_4000_4000_4000;
    #10 input_data = 256'h4200_4200_4200_4200_4200_4200_4200_42004200_4200_4200_42004200_4200_4200_4200;
    #10 input_data = 256'h4400_4400_4400_44004400_4400_4400_44004400_4400_4400_44004400_4400_4400_4400;
    #10input_data = 256'h3c00_3c00_3c00_3c00_3c00_3c00_3c00_3c003c00_3c00_3c00_3c003c00_3c00_3c00_3c00;
    #10 input_data = 0;
    #30 state = 1;
    
end

always begin
    #5 clk = ~clk;
end
    
endmodule
