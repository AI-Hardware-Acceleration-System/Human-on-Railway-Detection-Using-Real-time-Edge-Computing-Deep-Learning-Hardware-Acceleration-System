`timescale 1ns / 1ns
 
module PE16 #(parameter DATA_WIDTH = 16) (
    input logic clk,
    input logic rst_n,
    input logic [DATA_WIDTH-1:0] floatA,
    input logic [DATA_WIDTH-1:0] floatB,
    input logic [DATA_WIDTH-1:0] sum_in,
    output logic [DATA_WIDTH-1:0] sum_out
);

    logic [DATA_WIDTH-1:0] multResult;
    logic [DATA_WIDTH-1:0] addResult;    

    floatMult16 FM (
        .floatA(floatA),
        .floatB(floatB),
        .product(multResult)
    );

    floatAdd16 FADD (
        .floatA(multResult),
        .floatB(sum_in),
        .sum(addResult)
    );

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            //result_reg <= 0;
            sum_out <= 0;
        end else begin
            //result_reg <= result; // Store the previous value of result
            sum_out <= addResult;  // Update result
        end
    end
endmodule

module floatMult16 (
    input logic [15:0] floatA,
    input logic [15:0] floatB,
    output logic [15:0] product
);

    logic sign;
    logic signed [5:0] exponent; // 6th bit is the sign
    logic [9:0] mantissa;
    logic [10:0] fractionA, fractionB; // fraction = {1,mantissa}
    logic [21:0] fraction;

    always_comb begin
        if (floatA == 0 || floatB == 0) begin
            product = 0;
        end else begin
            sign = floatA[15] ^ floatB[15];
            exponent = floatA[14:10] + floatB[14:10] - 5'd15 + 5'd2;
        
            fractionA = {1'b1,floatA[9:0]};
            fractionB = {1'b1,floatB[9:0]};
            fraction = fractionA * fractionB;
            
            if (fraction[21] == 1'b1) begin
                fraction = fraction << 1;
                exponent = exponent - 1; 
            end else if (fraction[20] == 1'b1) begin
                fraction = fraction << 2;
                exponent = exponent - 2;
            end else if (fraction[19] == 1'b1) begin
                fraction = fraction << 3;
                exponent = exponent - 3;
            end else if (fraction[18] == 1'b1) begin
                fraction = fraction << 4;
                exponent = exponent - 4;
            end else if (fraction[17] == 1'b1) begin
                fraction = fraction << 5;
                exponent = exponent - 5;
            end else if (fraction[16] == 1'b1) begin
                fraction = fraction << 6;
                exponent = exponent - 6;
            end else if (fraction[15] == 1'b1) begin
                fraction = fraction << 7;
                exponent = exponent - 7;
            end else if (fraction[14] == 1'b1) begin
                fraction = fraction << 8;
                exponent = exponent - 8;
            end else if (fraction[13] == 1'b1) begin
                fraction = fraction << 9;
                exponent = exponent - 9;
            end else if (fraction[12] == 1'b0) begin
                fraction = fraction << 10;
                exponent = exponent - 10;
            end 
        
            mantissa = fraction[21:12];
            if(exponent[5]==1'b1) begin //exponent is negative
                product=16'b0000000000000000;
            end
            else begin
                product = {sign,exponent[4:0],mantissa};
            end
        end
    end
endmodule

module floatAdd16 (
    input logic [15:0] floatA,
    input logic [15:0] floatB,
    output logic [15:0] sum
);

    logic sign;
    logic signed [5:0] exponent; // 6th bit is the sign
    logic [9:0] mantissa;
    logic [4:0] exponentA, exponentB;
    logic [10:0] fractionA, fractionB, fraction; // fraction = {1,mantissa}
    logic [7:0] shiftAmount;
    logic cout;
    
    always_comb begin
        exponentA = floatA[14:10];
        exponentB = floatB[14:10];
        fractionA = {1'b1,floatA[9:0]};
        fractionB = {1'b1,floatB[9:0]}; 
        
        exponent = exponentA;
    
        if (floatA == 0) begin						//special case (floatA = 0)
            sum = floatB;
        end else if (floatB == 0) begin					//special case (floatB = 0)
            sum = floatA;
        end else if (floatA[14:0] == floatB[14:0] && floatA[15]^floatB[15]==1'b1) begin
            sum=0;
        end else begin
            if (exponentB > exponentA) begin
                shiftAmount = exponentB - exponentA;
                fractionA = fractionA >> (shiftAmount);
                exponent = exponentB;
            end else if (exponentA > exponentB) begin 
                shiftAmount = exponentA - exponentB;
                fractionB = fractionB >> (shiftAmount);
                exponent = exponentA;
            end
            if (floatA[15] == floatB[15]) begin			//same sign
                {cout,fraction} = fractionA + fractionB;
                if (cout == 1'b1) begin
                    {cout,fraction} = {cout,fraction} >> 1;
                    exponent = exponent + 1;
                end
                sign = floatA[15];
            end else begin						//different signs
                if (floatA[15] == 1'b1) begin
                    {cout,fraction} = fractionB - fractionA;
                end else begin
                    {cout,fraction} = fractionA - fractionB;
                end
                sign = cout;
                if (cout == 1'b1) begin
                    fraction = -fraction;
                end else begin
                end
                if (fraction [10] == 0) begin
                    if (fraction[9] == 1'b1) begin
                        fraction = fraction << 1;
                        exponent = exponent - 1;
                    end else if (fraction[8] == 1'b1) begin
                        fraction = fraction << 2;
                        exponent = exponent - 2;
                    end else if (fraction[7] == 1'b1) begin
                        fraction = fraction << 3;
                        exponent = exponent - 3;
                    end else if (fraction[6] == 1'b1) begin
                        fraction = fraction << 4;
                        exponent = exponent - 4;
                    end else if (fraction[5] == 1'b1) begin
                        fraction = fraction << 5;
                        exponent = exponent - 5;
                    end else if (fraction[4] == 1'b1) begin
                        fraction = fraction << 6;
                        exponent = exponent - 6;
                    end else if (fraction[3] == 1'b1) begin
                        fraction = fraction << 7;
                        exponent = exponent - 7;
                    end else if (fraction[2] == 1'b1) begin
                        fraction = fraction << 8;
                        exponent = exponent - 8;
                    end else if (fraction[1] == 1'b1) begin
                        fraction = fraction << 9;
                        exponent = exponent - 9;
                    end else if (fraction[0] == 1'b1) begin
                        fraction = fraction << 10;
                        exponent = exponent - 10;
                    end 
                end
            end
            mantissa = fraction[9:0];
            if(exponent[5]==1'b1) begin //exponent is negative
                sum = 16'b0000000000000000;
            end
            else begin
                sum = {sign,exponent[4:0],mantissa};
            end		
        end		
    end
endmodule

module adder_tree #(
    parameter int NUM_INPUTS = 8 // Number of inputs to the adder tree
) (
    input  logic [31:0] in[NUM_INPUTS],  // Array of 32-bit input numbers
    output logic [31:0] sum             // Final sum output
);

    // Determine the maximum number of stages required
    localparam int MAX_STAGES = $clog2(NUM_INPUTS);

    // Declare intermediate wires for each stage
    logic [31:0] stage_data[MAX_STAGES:0][NUM_INPUTS-1:0]; 

    // Stage 0: Assign initial inputs to stage_data
    initial begin
        for (int i = 0; i < NUM_INPUTS; i++) begin
            stage_data[0][i] = in[i];
        end
    end

    // Generate logic for each stage of the adder tree
    generate
        for (genvar stage = 0; stage < MAX_STAGES; stage++) begin
            for (genvar i = 0; i < (NUM_INPUTS >> (stage + 1)); i++) begin
                // Add pairs of numbers at the current stage
                always_comb stage_data[stage + 1][i] = 
                    stage_data[stage][2*i] + stage_data[stage][2*i + 1];
            end
            // Pass through remaining unpaired element, if any
            if ((NUM_INPUTS >> stage) % 2) begin
                always_comb stage_data[stage + 1][NUM_INPUTS >> (stage + 1)] = 
                    stage_data[stage][(NUM_INPUTS >> stage) - 1];
            end
        end
    endgenerate

    // Assign the final result
    assign sum = stage_data[MAX_STAGES][0];

endmodule

